magic
tech sky130A
magscale 1 2
timestamp 1717217591
<< pwell >>
rect 732 -382 794 -248
<< metal1 >>
rect 860 1314 1060 1406
rect 860 1310 1362 1314
rect 574 1250 1362 1310
rect 574 1246 1060 1250
rect 74 507 168 513
rect -468 -200 -268 -194
rect 74 -200 168 413
rect 320 134 384 140
rect -268 -400 200 -200
rect 320 -298 384 70
rect 320 -362 542 -298
rect -468 -406 -268 -400
rect 58 -574 198 -400
rect 574 -418 638 1246
rect 860 1206 1060 1246
rect 958 878 964 930
rect 1016 922 1022 930
rect 1016 886 1274 922
rect 1016 878 1022 886
rect 1148 750 1208 756
rect 935 507 1029 513
rect 935 333 1029 413
rect 962 286 1012 333
rect 681 236 1012 286
rect 681 -183 731 236
rect 1148 174 1208 690
rect 762 70 906 134
rect 970 70 976 134
rect 1092 114 1208 174
rect 762 -248 826 70
rect 1092 -186 1152 114
rect 732 -382 826 -248
rect 1168 -256 1190 -252
rect 1238 -256 1274 886
rect 854 -366 1080 -266
rect 1168 -358 1274 -256
rect 1302 -248 1362 1250
rect 2332 930 2384 936
rect 2332 872 2384 878
rect 1501 194 2076 195
rect 1490 64 2076 194
rect 1494 61 2076 64
rect 2210 61 2216 195
rect 1494 -190 1564 61
rect 2340 -180 2376 872
rect 2270 -204 2472 -180
rect 2270 -222 2830 -204
rect 2270 -240 2612 -222
rect 1302 -348 1508 -248
rect 1572 -336 2612 -240
rect 2768 -336 2830 -222
rect 1572 -346 2830 -336
rect 2270 -356 2830 -346
rect 1168 -362 1194 -358
rect 670 -574 730 -464
rect 58 -628 730 -574
rect 58 -1060 198 -628
rect 444 -806 644 -770
rect 854 -806 900 -366
rect 2270 -380 2472 -356
rect 1080 -770 1166 -460
rect 444 -902 900 -806
rect 986 -868 1186 -770
rect 444 -970 644 -902
rect 986 -928 1250 -868
rect 1310 -928 1368 -868
rect 986 -970 1186 -928
rect 1498 -1060 1576 -490
rect 58 -1194 1906 -1060
rect 66 -1198 1906 -1194
rect 2039 -1198 2045 -1060
<< via1 >>
rect 74 413 168 507
rect 320 70 384 134
rect -468 -400 -268 -200
rect 964 878 1016 930
rect 1148 690 1208 750
rect 935 413 1029 507
rect 906 70 970 134
rect 2332 878 2384 930
rect 2076 61 2210 195
rect 2612 -336 2768 -222
rect 1250 -928 1310 -868
rect 1906 -1198 2039 -1060
<< metal2 >>
rect 964 930 1016 936
rect 2326 922 2332 930
rect 1016 886 2332 922
rect 2326 878 2332 886
rect 2384 878 2390 930
rect 964 872 1016 878
rect -876 690 1148 750
rect 1208 690 1214 750
rect -876 -1288 -816 690
rect 68 413 74 507
rect 168 413 935 507
rect 1029 413 1035 507
rect 2076 195 2210 201
rect 906 134 970 140
rect 314 70 320 134
rect 384 70 906 134
rect 906 64 970 70
rect -474 -400 -468 -200
rect -268 -400 -262 -200
rect -468 -840 -268 -400
rect 1250 -868 1310 -862
rect 1310 -928 1368 -868
rect 1250 -934 1368 -928
rect -468 -1049 -268 -1040
rect 1308 -1288 1368 -934
rect 1906 -1060 2039 -1054
rect 2076 -1062 2210 61
rect 2814 -204 3259 -202
rect 2596 -222 3259 -204
rect 2596 -336 2612 -222
rect 2768 -336 3259 -222
rect 2596 -356 3259 -336
rect 3413 -356 3430 -202
rect 2039 -1195 2210 -1062
rect 1906 -1204 2039 -1198
rect -876 -1348 1368 -1288
<< via2 >>
rect -468 -1040 -268 -840
rect 3259 -356 3413 -202
<< metal3 >>
rect 3254 -202 3418 -197
rect 3254 -356 3259 -202
rect 3413 -319 4577 -202
rect 5373 -319 6247 -299
rect 3413 -356 6247 -319
rect 3254 -361 3418 -356
rect 4423 -600 6247 -356
rect -473 -840 -263 -835
rect -2520 -1040 -2514 -840
rect -2314 -1040 -468 -840
rect -268 -1040 -263 -840
rect 4423 -885 5550 -600
rect -473 -1045 -263 -1040
rect 4419 -1050 5550 -885
rect 6000 -1050 6247 -600
rect 4419 -1335 6247 -1050
<< via3 >>
rect -2514 -1040 -2314 -840
rect 5550 -1050 6000 -600
<< metal4 >>
rect 8057 -316 8893 -185
rect 5457 -327 6257 -319
rect 5363 -600 6257 -327
rect 8057 -600 8168 -316
rect -2515 -840 -2313 -839
rect -4884 -1040 -2514 -840
rect -2314 -1040 -2313 -840
rect -2515 -1041 -2313 -1040
rect 5363 -1050 5550 -600
rect 6000 -950 8168 -600
rect 8820 -950 8893 -316
rect 6000 -1050 8893 -950
rect 5363 -1317 6257 -1050
rect 8443 -1061 8893 -1050
<< via4 >>
rect -5204 -1100 -4884 -780
rect 8168 -950 8820 -316
<< metal5 >>
rect -28000 -780 -12000 7100
rect 15030 -128 31030 7066
rect 8046 -316 31030 -128
rect -5228 -780 -4860 -756
rect -28000 -1100 -5204 -780
rect -4884 -1100 -4860 -780
rect 8046 -950 8168 -316
rect 8820 -950 31030 -316
rect 8046 -1090 31030 -950
rect -28000 -9100 -12000 -1100
rect -5228 -1124 -4860 -1100
rect 15030 -9134 31030 -1090
<< glass >>
rect -27600 -8700 -12400 6700
rect 15430 -8734 30630 6666
use sky130_fd_pr__nfet_01v8_8HNZUS  XM1
timestamp 1717204734
transform 1 0 699 0 1 -324
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_5WKZCH  XM2
timestamp 1717204734
transform 1 0 1123 0 1 -328
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_J36GRF  XM3
timestamp 1717204734
transform 1 0 1537 0 1 -332
box -211 -310 211 310
<< labels >>
flabel metal1 2270 -380 2470 -180 0 FreeSans 256 0 0 0 VLow_Src
port 2 nsew
flabel metal1 444 -970 644 -770 0 FreeSans 256 0 0 0 VD_S
port 4 nsew
flabel metal1 860 1206 1060 1406 0 FreeSans 256 0 0 0 VD_H
port 0 nsew
flabel metal1 986 -970 1186 -770 0 FreeSans 256 0 0 0 VG_S
port 3 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 VG_H
port 1 nsew
<< end >>
